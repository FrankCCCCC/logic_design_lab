`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/29/2022 03:38:33 PM
// Design Name: 
// Module Name: segment7_frequency_divider
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`include "global.v"

//`define FREQ_DIV_BITS 30
// 1 Hz
//`define FREQ_DIV_COUNT `FREQ_DIV_BITS'd50000
//`define FREQ_DIV_COUNT `FREQ_DIV_BITS'd2
//`define FREQ_DIV_COUNT `FREQ_DIV_BITS'd5000000

module segment7_frequency_divider(
    clk_out,
    clk,
    rst
    );
    
    input clk;
    input rst;
    output clk_out;
    
    reg clk_in;
    reg clk_out;
    reg [`SEGMENT_7_FREQ_DIV_BITS-1:0] counter_in;
    reg [`SEGMENT_7_FREQ_DIV_BITS-1:0] counter_out;
    
    always@(counter_out or clk_out)
        if(counter_out < (`SEGMENT_7_FREQ_DIV_COUNT - 1))
        begin
            counter_in <= counter_out + `SEGMENT_7_FREQ_DIV_BITS'd1;
            clk_in <= clk_out;
        end
        else
        begin
            counter_in <= `SEGMENT_7_FREQ_DIV_BITS'd0;
            clk_in <= ~clk_out;
        end
        
    always@(posedge clk or negedge rst)
        if(~rst)
        begin
            counter_out <= `SEGMENT_7_FREQ_DIV_BITS'd0;
            clk_out <= 1'd0;
        end
        else
        begin
            counter_out <= counter_in;
            clk_out <= clk_in;
        end
endmodule
